`ifndef TEST_PKG_SVH
`define TEST_PKG_SVH

package test_pkg;

    `include "../../verification/tb/packet.sv"

    `include "../../verification/tb/cfg.sv"

    `include "../../verification/tb/gen.sv"

    `include "../../verification/tb/driver.sv"

    `include "../../verification/tb/monitor.sv"

    `include "../../verification/tb/agent.sv"

    `include "../../verification/tb/checker.sv"

    `include "../../verification/tb/env.sv"

    `include "../../verification/tb/test.sv"

endpackage

`endif  // TEST_PKG_SVH
