interface axis_uart_top_if;

bit clk_i;
bit arstn_i;

logic rx_i;
logic tx_o;

endinterface
