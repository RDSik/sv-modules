interface axil_if #(
    parameter int DATA_WIDTH = 32,
    parameter int ADDR_WIDTH = 32
) (
    input logic clk_i,
    input logic arstn_i
);

    localparam int STRB_WIDTH = (DATA_WIDTH / 8);

    logic [ADDR_WIDTH-1:0] awaddr;
    logic                  awvalid;
    logic                  awready;
    logic [           2:0] awprot;

    logic [DATA_WIDTH-1:0] wdata;
    logic [STRB_WIDTH-1:0] wstrb;
    logic                  wvalid;
    logic                  wready;

    logic [           1:0] bresp;
    logic                  bvalid;
    logic                  bready;

    logic [ADDR_WIDTH-1:0] araddr;
    logic                  arvalid;
    logic                  arready;
    logic [           2:0] arprot;

    logic [DATA_WIDTH-1:0] rdata;
    logic                  rvalid;
    logic                  rready;
    logic [           1:0] rresp;

    modport master(
        input clk_i,
        input arstn_i,
        output awaddr,
        output awprot,
        output awvalid,
        input awready,
        output wdata,
        output wstrb,
        output wvalid,
        input wready,
        input rresp,
        input bresp,
        input bvalid,
        output bready,
        output araddr,
        output arprot,
        output arvalid,
        input arready,
        input rdata,
        input rvalid,
        output rready
    );

    modport slave(
        input clk_i,
        input arstn_i,
        input awaddr,
        input awprot,
        input awvalid,
        output awready,
        input wdata,
        input wstrb,
        input wvalid,
        output wready,
        output rresp,
        output bresp,
        output bvalid,
        input bready,
        input araddr,
        input arprot,
        input arvalid,
        output arready,
        output rdata,
        output rvalid,
        input rready
    );

endinterface
