`ifndef TEST_PKG_SVH
`define TEST_PKG_SVH

package test_pkg;

    `include "packet.sv"

    `include "cfg.sv"

    `include "gen.sv"

    `include "driver.sv"

    `include "monitor.sv"

    `include "agent.sv"

    `include "checker.sv"

    `include "env.sv"

    `include "test.sv"

endpackage

`endif // TEST_PKG_SVH
