module axi_dma_wrap (
    axil_if.slave s_axil,

    axil_if.master m_axil_s2mm,
    axil_if.master m_axil_mm2s,

    axis_if.slave  s_axis_s2mm,
    axis_if.master m_axis_mm2s,

    output logic s2mm_introut_o,
    output logic mm2s_introut_o
);

    axi_dma_sim i_axi_dma_sim (
        .s_axi_lite_aclk       (s_axil.clk_i),
        .m_axi_mm2s_aclk       (m_axil_mm2s.clk_i),
        .m_axi_s2mm_aclk       (m_axil_s2mm.clk_i),
        .axi_resetn            (s_axil.arstn_i),
        .s_axi_lite_awvalid    (s_axil.awvalid),
        .s_axi_lite_awready    (s_axil.awready),
        .s_axi_lite_awaddr     (s_axil.awaddr),
        .s_axi_lite_wvalid     (s_axil.wvalid),
        .s_axi_lite_wready     (s_axil.wready),
        .s_axi_lite_wdata      (s_axil.wdata),
        .s_axi_lite_bresp      (s_axil.bresp),
        .s_axi_lite_bvalid     (s_axil.bvalid),
        .s_axi_lite_bready     (s_axil.bready),
        .s_axi_lite_arvalid    (s_axil.arvalid),
        .s_axi_lite_arready    (s_axil.arready),
        .s_axi_lite_araddr     (s_axil.araddr),
        .s_axi_lite_rvalid     (s_axil.rvalid),
        .s_axi_lite_rready     (s_axil.rready),
        .s_axi_lite_rdata      (s_axil.rdata),
        .s_axi_lite_rresp      (s_axil.rresp),
        .m_axi_mm2s_araddr     (m_axil_mm2s.araddr),
        .m_axi_mm2s_arlen      (),
        .m_axi_mm2s_arsize     (),
        .m_axi_mm2s_arburst    (),
        .m_axi_mm2s_arprot     (m_axil_mm2s.arprot),
        .m_axi_mm2s_arcache    (),
        .m_axi_mm2s_arvalid    (m_axil_mm2s.arvalid),
        .m_axi_mm2s_arready    (m_axil_mm2s.arready),
        .m_axi_mm2s_rdata      (m_axil_mm2s.rdata),
        .m_axi_mm2s_rresp      (m_axil_mm2s.rresp),
        .m_axi_mm2s_rlast      (),
        .m_axi_mm2s_rvalid     (m_axil_mm2s.rvalid),
        .m_axi_mm2s_rready     (m_axil_mm2s.rready),
        .mm2s_prmry_reset_out_n(),
        .m_axis_mm2s_tdata     (m_axis_mm2s.tdata),
        .m_axis_mm2s_tkeep     (m_axis_mm2s.tkeep),
        .m_axis_mm2s_tvalid    (m_axis_mm2s.tvalid),
        .m_axis_mm2s_tready    (m_axis_mm2s.tready),
        .m_axis_mm2s_tlast     (m_axis_mm2s.tlast),
        .m_axi_s2mm_awaddr     (m_axil_s2mm.awaddr),
        .m_axi_s2mm_awlen      (),
        .m_axi_s2mm_awsize     (),
        .m_axi_s2mm_awburst    (),
        .m_axi_s2mm_awprot     (m_axil_s2mm.awprot),
        .m_axi_s2mm_awcache    (),
        .m_axi_s2mm_awvalid    (m_axil_s2mm.awvalid),
        .m_axi_s2mm_awready    (m_axil_s2mm.awready),
        .m_axi_s2mm_wdata      (m_axil_s2mm.wdata),
        .m_axi_s2mm_wstrb      (m_axil_s2mm.wstrb),
        .m_axi_s2mm_wlast      (),
        .m_axi_s2mm_wvalid     (m_axil_s2mm.wvalid),
        .m_axi_s2mm_wready     (m_axil_s2mm.wready),
        .m_axi_s2mm_bresp      (m_axil_s2mm.bresp),
        .m_axi_s2mm_bvalid     (m_axil_s2mm.bvalid),
        .m_axi_s2mm_bready     (m_axil_s2mm.bready),
        .s2mm_prmry_reset_out_n(),
        .s_axis_s2mm_tdata     (s_axis_s2mm.tdata),
        .s_axis_s2mm_tkeep     (s_axis_s2mm.tkeep),
        .s_axis_s2mm_tvalid    (s_axis_s2mm.tvalid),
        .s_axis_s2mm_tready    (s_axis_s2mm.tready),
        .s_axis_s2mm_tlast     (s_axis_s2mm.tlast),
        .mm2s_introut          (mm2s_introut_o),
        .s2mm_introut          (s2mm_introut_o),
        .axi_dma_tstvec        ()
    );

endmodule
