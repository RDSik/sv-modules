`timescale 1ns / 1ps

`include "modules/spi/tb/axil_spi_class.svh"
`include "modules/uart/tb/axil_uart_class.svh"
`include "modules/i2c/tb/axil_i2c_class.svh"
`include "modules/rgmii/tb/axil_rgmii_class.svh"

module axil_top_tb ();

    localparam int FIFO_DEPTH = 128;
    localparam int CS_WIDTH = 8;
    localparam int RGMII_WIDTH = 4;
    localparam int AXIL_ADDR_WIDTH = 32;
    localparam int AXIL_DATA_WIDTH = 32;
    localparam int AXIS_DATA_WIDTH = 8;
    localparam int MASTER_NUM = 1;
    localparam int SLAVE_NUM = 4;

    localparam logic [AXIL_ADDR_WIDTH-1:0] BASE_LOW_ADDR = 32'h43c0_0000;
    localparam logic [AXIL_ADDR_WIDTH-1:0] BASE_HIGTH_ADDR = 32'h43c0_ffff;
    localparam logic [AXIL_ADDR_WIDTH-1:0] ADDR_OFFSET = 32'h0001_0000;

    function automatic logic [SLAVE_NUM-1:0][AXIL_ADDR_WIDTH-1:0] slave_addr_get;
        input logic [AXIL_ADDR_WIDTH-1:0] addr;
        begin
            for (int i = 0; i < SLAVE_NUM; i++) begin
                slave_addr_get[i] = addr + i * ADDR_OFFSET;
            end
        end
    endfunction

    localparam logic [SLAVE_NUM-1:0][AXIL_ADDR_WIDTH-1:0] SLAVE_LOW_ADDR = slave_addr_get(
        BASE_LOW_ADDR
    );
    localparam logic [SLAVE_NUM-1:0][AXIL_ADDR_WIDTH-1:0] SLAVE_HIGH_ADDR = slave_addr_get(
        BASE_HIGTH_ADDR
    );

    localparam int WAT_CYCLES = 250;
    localparam int CLK_PER_NS = 2;
    localparam int RESET_DELAY = 10;

    logic clk_i;
    logic arstn_i;
    logic uart;

    spi_if #(.CS_WIDTH(CS_WIDTH)) m_spi ();

    assign m_spi.miso = m_spi.mosi;

    eth_if #(.DATA_WIDTH(RGMII_WIDTH)) m_eth ();

    assign m_eth.rxd    = m_eth.txd;
    assign m_eth.rx_ctl = m_eth.tx_ctl;
    assign m_eth.rx_clk = clk_i;

    axis_if #(
        .DATA_WIDTH(AXIS_DATA_WIDTH)
    ) m_axis (
        .clk_i(clk_i),
        .rst_i(~arstn_i)
    );

    axis_if #(
        .DATA_WIDTH(AXIS_DATA_WIDTH)
    ) s_axis (
        .clk_i(clk_i),
        .rst_i(~arstn_i)
    );

    axil_if #(
        .ADDR_WIDTH(AXIL_ADDR_WIDTH),
        .DATA_WIDTH(AXIL_DATA_WIDTH)
    ) s_axil[MASTER_NUM-1:0] (
        .clk_i  (clk_i),
        .arstn_i(arstn_i)
    );

    initial begin
        arstn_i = 1'b0;
        repeat (RESET_DELAY) @(posedge clk_i);
        arstn_i = 1'b1;
        $display("Reset done in: %0t ns\n.", $time());
    end

    initial begin
        clk_i = 1'b0;
        forever begin
            #(CLK_PER_NS / 2) clk_i = ~clk_i;
        end
    end

    initial begin
        axil_uart_class #(
            .DATA_WIDTH(AXIL_DATA_WIDTH),
            .ADDR_WIDTH(AXIL_ADDR_WIDTH),
            .BASE_ADDR (SLAVE_LOW_ADDR[0])
        ) uart;
        axil_spi_class #(
            .DATA_WIDTH(AXIL_DATA_WIDTH),
            .ADDR_WIDTH(AXIL_ADDR_WIDTH),
            .BASE_ADDR (SLAVE_LOW_ADDR[1])
        ) spi;
        axil_i2c_class #(
            .DATA_WIDTH(AXIL_DATA_WIDTH),
            .ADDR_WIDTH(AXIL_ADDR_WIDTH),
            .BASE_ADDR (SLAVE_LOW_ADDR[2])
        ) i2c;
        axil_rgmii_class #(
            .DATA_WIDTH(AXIL_DATA_WIDTH),
            .ADDR_WIDTH(AXIL_ADDR_WIDTH),
            .TLAST_EN  (0),
            .BASE_ADDR (SLAVE_LOW_ADDR[3])
        ) rgmii;
        uart  = new(s_axil[0]);
        spi   = new(s_axil[0]);
        rgmii = new(s_axil[0], m_axis, s_axis);
        i2c   = new(s_axil[0]);
        uart.uart_start();
        spi.spi_start();
        i2c.i2c_start();
        rgmii.rgmii_start();
        $stop;
    end

    initial begin
        $dumpfile("axil_top_tb.vcd");
        $dumpvars(0, axil_top_tb);
    end

    axil_top #(
        .AXIL_ADDR_WIDTH(AXIL_ADDR_WIDTH),
        .AXIL_DATA_WIDTH(AXIL_DATA_WIDTH),
        .FIFO_DEPTH     (FIFO_DEPTH),
        .SPI_CS_WIDTH   (CS_WIDTH),
        .RGMII_WIDTH    (RGMII_WIDTH),
        .SLAVE_NUM      (SLAVE_NUM),
        .MASTER_NUM     (MASTER_NUM),
        .SLAVE_LOW_ADDR (SLAVE_LOW_ADDR),
        .SLAVE_HIGH_ADDR(SLAVE_HIGH_ADDR),
        .ILA_EN         (0),
        .MODE           ("sync"),
        .VENDOR         ("")
    ) i_axil_top (
        .clk_i    (clk_i),
        .uart_rx_i(uart),
        .uart_tx_o(uart),
        .s_axil   (s_axil),
        .s_axis   (m_axis),
        .m_axis   (s_axis),
        .m_spi    (m_spi),
        .m_eth    (m_eth)
    );

endmodule
