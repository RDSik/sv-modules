/* verilator lint_off TIMESCALEMOD */
module fir_filter #(
    parameter     COE_FILE   = "fir.mem",
    parameter int CH_NUM     = 2,
    parameter int DATA_WIDTH = 16,
    parameter int COEF_WIDTH = 18,
    parameter int TAP_NUM    = 4
) (
    input logic clk_i,
    input logic rstn_i,
    input logic en_i,

    input logic                                     tvalid_i,
    input logic signed [CH_NUM-1:0][DATA_WIDTH-1:0] tdata_i,

    output logic                                                        tvalid_o,
    output logic signed [CH_NUM-1:0][COEF_WIDTH+DATA_WIDTH+TAP_NUM-1:0] tdata_o
);

    logic [COEF_WIDTH-1:0] coe_mem[TAP_NUM];

    initial begin
        $readmemh(COE_FILE, coe_mem);
    end

    localparam int DELAY = 2 * TAP_NUM;

    logic [DELAY-1:0] tvalid_d;

    always_ff @(posedge clk_i) begin
        if (~rstn_i) begin
            tvalid_d <= '0;
        end else begin
            tvalid_d <= {tvalid_d[DELAY-2:0], tvalid_i};
        end
    end

    always_ff @(posedge clk_i) begin
        if (~rstn_i) begin
            tvalid_o <= 1'b0;
        end else begin
            if (en_i) begin
                tvalid_o <= tvalid_d[DELAY-1];
            end else begin
                tvalid_o <= 1'b0;
            end
        end
    end

    for (genvar ch_indx = 0; ch_indx < CH_NUM; ch_indx++) begin : g_ch
        logic signed [TAP_NUM-1:0][                   DATA_WIDTH-1:0] delay;
        logic signed [TAP_NUM-1:0][        DATA_WIDTH+COEF_WIDTH-1:0] mult;
        logic signed [TAP_NUM-1:0][DATA_WIDTH+COEF_WIDTH+TAP_NUM-1:0] acc;

        always_ff @(posedge clk_i) begin
            if (tvalid_i) begin
                delay[0] <= tdata_i[ch_indx];
            end
            for (int tap_indx = 1; tap_indx < TAP_NUM; tap_indx++) begin
                delay[tap_indx] <= delay[tap_indx-1];
            end
        end

        always_ff @(posedge clk_i) begin
            for (int tap_indx = 0; tap_indx < TAP_NUM; tap_indx++) begin
                mult[tap_indx] <= delay[tap_indx] * coe_mem[tap_indx];
            end
        end

        always_ff @(posedge clk_i) begin
            acc[0] <= mult[0];
            for (int tap_indx = 1; tap_indx < TAP_NUM; tap_indx++) begin
                acc[tap_indx] <= mult[tap_indx] + acc[tap_indx-1];
            end
        end

        always_ff @(posedge clk_i) begin
            tdata_o[ch_indx] <= acc[TAP_NUM-1];
        end
    end

endmodule
