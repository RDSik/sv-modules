`ifndef TEST_PKG_SVH
`define TEST_PKG_SVH

package test_pkg;
    `include "../../verification/tb/cfg.svh"
    `include "../../verification/tb/env.svh"
endpackage

`endif  // TEST_PKG_SVH
