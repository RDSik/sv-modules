interface axis_uart_top_if;

bit clk_i;
bit arstn_i;

logic uart_rx_i;
logic uart_tx_o;

endinterface
