`ifndef PACKET_SV
`define PACKET_SV

class packet;
    rand logic [7:0] tdata;
    rand int         delay;
endclass

`endif // PACKET_SV
